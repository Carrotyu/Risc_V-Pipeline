module Instruction_Memory(rst, clk, read_address, instruction_out);

input rst, clk;
input [31:0] read_address;
output [31:0] instruction_out;
reg [31:0] I_Mem [63:0];  
integer k;
assign instruction_out = I_Mem[read_address];

always @(posedge clk or posedge rst)
begin
    if (rst) begin
        for (k = 0; k < 64; k = k + 1) begin 
            I_Mem[k] = 32'b00;  
        end
    end else begin
        // R-type
        I_Mem[0] = 32'b0000000000000000000000000000000 ;       // no operation
        I_Mem[4] = 32'b00000001100110000000011010110011;    // add x13, x16, x25
        I_Mem[8] = 32'b01000000001101000000001010110011;     // sub x5, x8, x3
        I_Mem[12] = 32'b00000000001100010111000010110011;    // and x1, x2, x3
        I_Mem[16] = 32'b00000000010100011110001000110011;    // or x4, x3, x5
        I_Mem[20] = 32'b00000000010100011100001000110011;    // xor x4, x3, x5
	I_Mem[24] = 32'b00000000010100011001001000110011;    // sll x4, x3, x5
        I_Mem[28] = 32'b00000000010100011101001000110011;    // srl x4, x3, x5
        I_Mem[32] = 32'b01000000001000011101001010110011;    //sra x5, x3, x2
        I_Mem[36] = 32'b00000000001000011010001010110011;    //slt x5, x3, x2 
        // I-type
        I_Mem[40]  = 32'b00000000001010101000101100010011;     // addi x22, x21, 2
        I_Mem[44]  = 32'b00000000001101000110010010010011;     // ori x9, x8, 3 
	I_Mem[48] = 32'b00000000010001000110010010010011;     // xori x9, x8, 4
	I_Mem[52] = 32'b00000000010100010111000010010011;     // andi x1, x2, 5
	I_Mem[56] = 32'b00000000011000011001001000010011;    // slli x4, x3, 6
	I_Mem[60] = 32'b00000000011100011101001000010011;    // srli x4, x3, 7 
	I_Mem[64] = 32'b00000000100000011101001010010011;    //srai x5, x3, 8
	I_Mem[68] = 32'b00000000100100011010001010010011;    //slti x5, x3, 9  
        // L-type
	I_Mem[72]=  32'b00000000010100011000010010000011;     // lb x9, 5(x3)
	I_Mem[76] = 32'b00000000001100011001010010000011;    // lh x9, 3(x3)
        I_Mem[80]= 32'b00000000111100010010010000000011;    // lw x8, 15(x2) 
        // S-type
        I_Mem[84] =  32'b00000000111100011000010000100011;     // sb x15, 8(x3), x3 = 12
	I_Mem[86] =  32'b00000000111000110001010100100011;     // sh x14, 10(x6), x6 = 44
	I_Mem[90] = 32'b00000000111000110010011000100011;     // sw x14, 12(x6), x6 = 44     
	//B-type    
	I_Mem[94] = 32'b00000000100101001000011001100011;     // beq x9, x9, 12, (PC + 12 if x9 = x9 
	I_Mem[98] = 32'b00000000100101001001011101100011;     //bne x9, x9, 14,(PC + 14 if x9 != x9)
	// U-type
        I_Mem[102] =  32'b00000000000000101000000110110111;     // lui x3, 40
        I_Mem[106] =  32'b0000000000000010100001010010111;     // auipc x5, 20 (rd = PC + (imm << 12))
	// J-type
	I_Mem[110] = 32'b0_0000000000000010100_000011101111;         // jal x1, 20


        
    end
end

endmodule
